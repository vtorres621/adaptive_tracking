b0VIM 8.1      �fa�A �  root                                    xilinx-zcu102-2020_2                    ~root/eco/pytracking/tracker/eco/eco.py                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            3210    #"! U                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 tp           V                            M       W              	       Q       �                            �                     E                           V       R                    V       �                           �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     ad  C   �     V       �  �  �  �  ^  &  �  �  �  J    
  �  �  �  �  �  �  �  �  c  5      
  �  �  �  q  p  P  5    �  �  �  f  H  %  $    �
  �
  �
  R
  Q
  1
  �	  �	  �	  ~	  ^	  	  �  n  0  �  �  �  n  m  :  �  w      �  �  n  )  �  l  k  O         �  �  w    �      �  �  �                                                                             #print("[INFO][eco.py] get regularization filter")         # Get regularization filter                                                  self.params.interpolation_windowing, self.params.device) for sz in self.filter_sz])                                                 self.params.interpolation_bicubic_a, self.params.interpolation_centering,         self.interp_fs = TensorList([dcf.get_interp_fourier(sz, self.params.interpolation_method,         # Get interpolation function          self.window = TensorList([dcf.hann2d(sz).to(self.params.device) for sz in self.feature_sz])         # Get window function          self.num_filters = len(self.filter_sz)         # Number of filters          self.compressed_dim = self.fparams.attribute('compressed_dim')         self.output_sz = self.params.score_upsample_factor * self.img_support_sz    # Interpolated size of the output         self.filter_sz = self.feature_sz + (self.feature_sz + 1) % 2         self.feature_sz = self.params.features.size(self.img_sample_sz)         self.img_support_sz = self.img_sample_sz         # Set other sizes (corresponds to ECO code)          self.img_sample_sz += feat_max_stride - self.img_sample_sz % (2 * feat_max_stride)         self.img_sample_sz = torch.round(torch.sqrt(torch.prod(self.base_target_sz * self.params.search_area_scale))) * torch.ones(2)         feat_max_stride = max(self.params.features.stride())         # Use odd square search area and set sizes          self.base_target_sz = self.target_sz / self.target_scale         # Target size in base scale              self.target_scale =  math.sqrt(search_area / self.params.min_image_sample_size)         elif search_area < self.params.min_image_sample_size:             self.target_scale =  math.sqrt(search_area / self.params.max_image_sample_size)         if search_area > self.params.max_image_sample_size:         search_area = torch.prod(self.target_sz * self.params.search_area_scale).item()         self.target_scale = 1.0         # Set search area          self.target_sz = torch.Tensor([state[3], state[2]])         self.pos = torch.Tensor([state[1] + (state[3] - 1)/2, state[0] + (state[2] - 1)/2])         # Get position and size          self.fparams = self.params.features.get_fparams('feature_params')         # Get feature specific params          self.params.features.set_is_color(image.shape[2] == 3)         # Chack if image is color          self.initialize_features()         # Initialize features         #print(self.params.device)             self.params.device = 'cpu' if self.params.use_gpu else 'cpu'         if not self.params.has('device'):         #print("THERE")         #self.params.use_gpu = 0         self.frame_num = 1         # Initialize some stuff          state = info['init_bbox']          #print("[INFO][eco.py] initialize called")     def initialize(self, image, info: dict, dpu_features) -> dict:           self.features_initialized = True             self.params.features.initialize()         if not getattr(self, 'features_initialized', False):     def initialize_features(self):      multiobj_mode = 'parallel'  class ECO(BaseTracker):   import time import numpy as np from pytracking.features import augmentation from .optim import FilterOptim, FactorizedConvProblem from pytracking.libs.optimization import GaussNewtonCG from pytracking.utils.plotting import show_tensor from pytracking.features.preprocessing import numpy_to_torch from pytracking.libs.tensorlist import tensor_operation from pytracking import complex, dcf, fourier, TensorList import math import torch.nn.functional as F import torch from pytracking.tracker.base import BaseTracker ad  y  �            �  �  �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       hf[:,:,:,0,:] += complex.conj(hf[:,:,:,0,:].flip((2,)))             hf[:,:,:,0,:] /= 2 ad  �  
            �  �  �       �  �  �  �  �  n  m  G  �  �  �  �  �  N  M  
  	    �  L  
    A    �  �  �  �  �  �  D  �
  �
  
  ~
  }
  Z
  Y
  X
  =
  �	  �	  �	  �	  �	  Z	  	  	  	   	  �  �  �  �  �  @        �  �  f  e  <  �  �  �  �  �  �  >  =    �  �  K  	  �  v  ;  �  �  ~  K    �  �  �  $  �                                                                                              (math.floor(pd[1].item()), math.ceil(pd[1].item()),                     scores_scales.append(F.pad(fourier.sample_fs(sfe[sind:sind+1,...], sz),                     pd = (self.output_sz-sz)/2                 for sind, sz in enumerate(sample_sz):                 scores_scales = []                 sfe = fourier.shift_fs(sfe, math.pi*torch.ones(2))             for sfe, a, b in zip(sf, alpha, beta):             scores = 0             sample_sz = torch.round(self.output_sz.view(1,-1) * self.params.scale_factors.view(-1,1))             beta = self.fparams.attribute('translation_weight')             alpha = self.fparams.attribute('scale_weight')         elif self.params.score_fusion_strategy == 'transcale':             scores = fourier.sample_fs(fourier.sum_fs(weight * sf), self.output_sz)             weight = self.fparams.attribute('translation_weight')         elif self.params.score_fusion_strategy == 'weightedsum':             scores = fourier.sample_fs(fourier.sum_fs(sf), self.output_sz)         if self.params.score_fusion_strategy == 'sum':     def localize_target(self, sf: TensorList):          return complex.mult(self.filter, sample_xf).sum(1, keepdim=True)     def apply_filter(self, sample_xf: TensorList) -> torch.Tensor:           return out, sample_pos, sample_scales          #print("[TIME][eco.py] Track end: ", track_end - track4)         #track_end = time.perf_counter()          out = {'target_bbox': new_state.tolist()}         new_state = torch.cat((self.pos[[1,0]] - (self.target_sz[[1,0]]-1)/2, self.target_sz[[1,0]]))         # Return new state               self.symmetrize_filter()             self.filter_optimizer.run(self.params.CG_iter, train_xf)         if self.frame_num % self.params.train_skipping == 1:         # Train filter           self.update_memory(train_xf)         # Update memory           train_xf = fourier.shift_fs(train_xf, shift=shift_samp)         shift_samp = 2*math.pi * (self.pos - sample_pos) / (sample_scales[scale_ind] * self.img_support_sz)         # Shift the sample                   train_xf = TensorList([xf[scale_ind:scale_ind+1, ...] for xf in test_xf])         # Get train sample           # ------- UPDATE ------- #               show_tensor(score_map, 5, title='Max score = {:.2f}'.format(max_score))         elif self.params.debug >= 2:             self.visdom.register(self.debug_info, 'info_dict', 1, 'Status')             self.visdom.register(score_map, 'heatmap', 2, 'Score Map')         if self.visdom is not None:                    self.debug_info['max_score'] = max_score         max_score = torch.ma           print("[INFO][eco.py][track] Pos_updated: ", pos_updated)         pos_updated, target_scale_updated, target_sz_updated = self.update_state(sample_pos + translation_vec, self.target_scale * scale_change_factor)         # Update position and scale           scale_change_factor = self.params.scale_factors[scale_ind]          #print("[TIME][eco.py][track] Checkpoint 4: ", track4 - track3)         #track4 = time.perf_counter()          translation_vec, scale_ind, s = self.localize_target(sf)          #print("[TIME][eco.py][track] Checkpoint 3: ", track3 - track2)         #track3 = time.perf_counter()          sf = self.apply_filter(test_xf)         # Compute scores           #print("[TIME][eco.py][track] Checkpoint 2: ", track2 - track1)         #track2 = time.perf_counter()          test_xf = self.extract_fourier_sample(dpu_features,im, self.pos, sample_scales, self.img_sample_sz)          #print("[TIME][eco.py][track] Checkpoint 1: ", track1 - track_start)         #track1 = time.perf_counter() ad  U  �     E       �  �  �  �  w  n  m  l  H    �  �  <  ;  :        �  �  �  �  �  �    �  �  �  �  �  �  �    B  �  �  �  �  �  U  #  "  �
  �
  �
  �
  �
  �
  D
  �	  �	  �	  �	  I	  	  �  r  3  �  �  R  ;    �  �  l  =  �  �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   (math.floor(pd[1].item()), math.ceil(pd[1].item()),                     scores_scales.append(F.pad(fourier.sample_fs(sfe[sind:sind+1,...], sz),                     pd = (self.output_sz-sz)/2                 for sind, sz in enumerate(sample_sz):                 scores_scales = []                 sfe = fourier.shift_fs(sfe, math.pi*torch.ones(2))             for sfe, a, b in zip(sf, alpha, beta):             scores = 0             sample_sz = torch.round(self.output_sz.view(1,-1) * self.params.scale_factors.view(-1,1))             beta = self.fparams.attribute('translation_weight')             alpha = self.fparams.attribute('scale_weight')         elif self.params.score_fusion_strategy == 'transcale':             scores = fourier.sample_fs(fourier.sum_fs(weight * sf), self.output_sz)             weight = self.fparams.attribute('translation_weight')         elif self.params.score_fusion_strategy == 'weightedsum':             scores = fourier.sample_fs(fourier.sum_fs(sf), self.output_sz)         if self.params.score_fusion_strategy == 'sum':     def localize_target(self, sf: TensorList):          return complex.mult(self.filter, sample_xf).sum(1, keepdim=True)     def apply_filter(self, sample_xf: TensorList) -> torch.Tensor:           return out, sample_pos, sample_scales          #print("[TIME][eco.py] Track end: ", track_end - track4)         #track_end = time.perf_counter()          out = {'target_bbox': new_state.tolist()}         new_state = torch.cat((self.pos[[1,0]] - (self.target_sz[[1,0]]-1)/2, self.target_sz[[1,0]]))         # Return new state               self.symmetrize_filter()             self.filter_optimizer.run(self.params.CG_iter, train_xf)         if self.frame_num % self.params.train_skipping == 1:         # Train filter           self.update_memory(train_xf)         # Update memory           train_xf = fourier.shift_fs(train_xf, shift=shift_samp)         shift_samp = 2*math.pi * (self.pos - sample_pos) / (sample_scales[scale_ind] * self.img_support_sz)         # Shift the sample                   train_xf = TensorList([xf[scale_ind:scale_ind+1, ...] for xf in test_xf])         # Get train sample           # ------- UPDATE ------- #               show_tensor(score_map, 5, title='Max score = {:.2f}'.format(max_score))         elif self.params.debug >= 2:             self.visdom.register(self.debug_info, 'info_dict', 1, 'Status')             self.visdom.register(score_map, 'heatmap', 2, 'Score Map')         if self.visdom is not None:                    self.debug_info['max_score'] = max_score         max_score = torch.max(score_map).item()         score_map = s[scale_ind, ...]   ad  &   �     V       �  l  
  �  �  �  �  v  C      �  �  B    �  �  �    �  �  �  `  _  ^  �
  �
  �
  "
  !
  �	  �	  �	  �	  �	  H	  G	  $	  #	  �  �  �  �  �  f  !             �  �  �  Q    �  �  ~  Y    �  }  |  O  5  �  �  �  �  �  b  ,  +  �  �  �  �  N  /     �  `    �  �  �                                                if 'rotate' in self.params.augmentation:             transforms.append(augmentation.FlipHorizontal())         if 'fliplr' in self.params.augmentation and self.params.augmentation['fliplr']:             transforms.extend([augmentation.Translation(shift) for shift in self.params.augmentation['shift']])         if 'shift' in self.params.augmentation:         transforms = [augmentation.Identity()]         # Do data augmentation     def generate_init_samples(self, im: torch.Tensor, dpu_features) -> TensorList:          return _project_sample(x, self.projection_matrix)              return torch.matmul(x.permute(2, 3, 0, 1), P).permute(2, 3, 0, 1)              #print("[INFO][eco.py] x:\n", x[0][0][0])             #print("[INFO][eco.py] P:\n", P)                  return x                 #print("[INFO][eco.py] P is None")             if P is None:         def _project_sample(x: torch.Tensor, P: torch.Tensor):         @tensor_operation     def project_sample(self, x: TensorList):          return TensorList([dcf.interpolate_dft(xf, bf) for xf, bf in zip(sample_xf, self.interp_fs)])         #np.save('hw_samplexf', sample_xf[0][0][0])         #print("[INFO][eco.py] sample_xf:\n", sample_xf[0][0][0])         sample_xf = fourier.cfft2(x)         #np.save('hw_x*window', x[0][0][0])         #print("[INFO][eco.py] x *= self. window:\n", x[0][0][0][0])         x *= self.window         #print("[INFO][eco.py] self.window:\n", self.window[0][0][0][0])         #print("[INFO][eco.py] x:\n", x[0][0][0][0])     def preprocess_sample(self, x: TensorList) -> TensorList:          #return self.preprocess_sample(self.project_sample(x))         return x                     #print("[TIME][eco.py][fourier] CP1: ", fourier4 - fourier3)         #fourier4 = time.perf_counter()          x = self.preprocess_sample(x)          #print("[TIME][eco.py][fourier] CP1: ", fourier3 - fourier2)         #fourier3 = time.perf_counter()          x = self.project_sample(x)          #print("[TIME][eco.py][fourier] CP1: ", fourier2 - fourier1)         #fourier2 = time.perf_counter()          x = self.extract_sample(dpu_features,im, pos, scales, sz)          #fourier1 = time.perf_counter()      def extract_fourier_sample(self, dpu_features,im: torch.Tensor, pos: torch.Tensor, scales, sz: torch.Tensor) -> TensorList:          return self.params.features.extract(dpu_features,im, pos, scales, sz)[0]     def extract_sample(self, dpu_features,im: torch.Tensor, pos: torch.Tensor, scales, sz: torch.Tensor):           return translation_vec, scale_ind, scores              translation_vec *= self.params.scale_factors[scale_ind]         if self.params.score_fusion_strategy in ['sum', 'weightedsum']:         translation_vec = disp[scale_ind, ...].view(-1) * (self.img_support_sz / self.output_sz) * self.target_scale         # Compute translation vector and scale change factor              disp = max_disp - self.output_sz / 2         elif self.params.score_fusion_strategy == 'transcale':             disp = (max_disp + self.output_sz / 2) % self.output_sz - self.output_sz / 2         if self.params.score_fusion_strategy in ['sum', 'weightedsum']:         # Convert to displacements in the base scale          max_disp = max_disp.float().cpu()         _, scale_ind = torch.max(max_score, dim=0)         max_score, max_disp = dcf.max2d(scores)         # Get maximum              raise ValueError('Unknown score fusion strategy.')         else:                 scores = scores + (b - a) * scores_cat.mean(dim=0, keepdim=True) + a * scores_cat                 scores_cat = torch.cat(scores_scales)                                          math.floor(pd[0].item()), math.ceil(pd[0].item())))) ad      �     V       �  e  �  �  �  ~  }  �  �  �  h  g  b  9    �  �  ^  B    �  �  f  Y    �
  �
  �
  
  �	  �	  �	  �	  �	  �	  	  M	  	  �  }  |  {  V  =  �  v  \  B  (    �  �  �  �  |  W  #  �  �  �  �  p  J  I    �  �  �  �  ^  G  �  �  �  �  {  =  �  �  �  c    �  �  �  �  �                                          for hf in self.filter:     def symmetrize_filter(self):          return pos_updated, target_scale_updated, target_sz_updated         #print("[INFO][eco.py] update_state pos_updated:\n", pos_updated)         target_sz_updated = self.target_sz         target_scale_updated = self.target_scale         pos_updated = self.pos         self.pos = torch.max(torch.min(new_pos, self.image_sz - inside_offset), inside_offset)         inside_offset = (inside_ratio - 0.5) * self.target_sz         inside_ratio = 0.2         # Update pos          self.target_sz = self.base_target_sz * self.target_scale         self.target_scale = new_scale.clamp(self.min_scale_factor, self.max_scale_factor)         # Update scale         #print("[INFO][eco.py] update_state new_pos: \n", new_pos)     def update_state(self, new_pos, new_scale):          return replace_ind         self.num_stored_samples += 1         self.previous_replace_ind = replace_ind.copy()              replace_ind.append(r_ind)             sw /= sw.sum()                      sw[r_ind] = sw[prev_ind] / (1 - fparams.learning_rate)                 else:                     sw[r_ind] = fparams.learning_rate                     sw /= 1 - fparams.learning_rate                 if prev_ind is None:                 # Update weights                  r_ind = r_ind.item()                 _, r_ind = torch.min(sw, 0)                 # Get index to replace             else:                 r_ind = 0                 sw[0] = 1                 sw[:] = 0             if num_samp == 0 or fparams.learning_rate == 1:         for sw, prev_ind, num_samp, fparams in zip(self.sample_weights, self.previous_replace_ind, self.num_stored_samples, self.fparams):         replace_ind = []     def update_sample_weights(self):               train_samp[:,:,ind:ind+1,:,:] = xf.permute(2, 3, 0, 1, 4)         for train_samp, xf, ind in zip(self.training_samples, sample_xf, replace_ind):         replace_ind = self.update_sample_weights()         # Update weights and get index to replace     def update_memory(self, sample_xf: TensorList):           return init_samples           #np.save('hw_init_samples2', init_samples[0][0][0])                     init_samples[i] = torch.cat([init_samples[i], F.dropout2d(init_samples[i][0:1,...].expand(num,-1,-1,-1), p=prob, training=True)])                     #print(init_samples[i].shape)                 if use_aug:                              for i, use_aug in enumerate(self.fparams.attribute('use_augmentation')):                          num, prob = self.params.augmentation['dropout']         if 'dropout' in self.params.augmentation:         #print("DONE REMOVING AUGMENTED SAMPLES")                 init_samples[i] = init_samples[i][0:1, ...]             if not use_aug:         for i, use_aug in enumerate(self.fparams.attribute('use_augmentation')):         # Remove augmented samples for those that shall not have         #print(init_samples.size)         #print("SIZE OF INIT_SAMPLES")         #init_samples = ([dpu_features])               #np.save('hw_init_samples1', init_samples[0][0][0])         #print("[INFO][eco.py] init_samples: \n", init_samples[0][0][0])          init_samples = self.params.features.extract_transformed(im, self.pos, self.target_scale, self.img_sample_sz, transforms, dpu_features)          #print("[INFO][eco.py] self.target_scale: ", self.target_scale)         #print("[INFO][eco.py] self.pos: ", self.pos)              transforms.extend([augmentation.Blur(sigma) for sigma in self.params.augmentation['blur']])         if 'blur' in self.params.augmentation:             transforms.extend([augmentation.Rotate(angle) for angle in self.params.augmentation['rotate']]) ad  -   }     M       }  9  8  �  �  �  �  
  �  �  m    �  �  u  �  �  �  �  �  �  �  `    �
  �
  �
  n
  6
  �	  �	  �	  �	  �	  u	  	  �  �  �  `  W  &  �  �  �  �  �  p  g  f  5  ,  �  N  �  �  b    �  �  �  p  "  �  �  ^  "  �  �  �  �  �  f  A  $  �  }  |                                                                   shift_samp = 2 * math.pi * torch.Tensor(shift) / self.img_support_sz                 for i, shift in enumerate(self.params.augmentation['shift']):                     continue                 if xf.shape[0] == 1:             for xf in train_xf:         if 'shift' in self.params.augmentation:         # Shift the samples back                  #brea         #np.save('hw_train_xf1', train_xf[1][0][0])         #print("[INFO][eco.py] train_xf[1]: ", train_xf[1])         #print("[INFO][eco.py] train_xf[1] shape: ", train_xf[1][0][0].shape)         #np.save('hw_train_xf0', train_xf[0][0][0])         #print("[INFO][eco.py] train_xf[0]: ", train_xf[0].shape)         #print("[INFO][eco.py] train_xf[0] shape: ", train_xf[0][0][0].shape)         train_xf = self.preprocess_sample(x)         # Transform to get the training sample                  #np.save('hw_proj1', self.projection_matrix[1])         #print("[INFO][eco.py] projection matrix[1]: \n", self.projection_matrix[1])         #print("[INFO][eco.py] projection matrix[1]shape : ", self.projection_matrix[1].shape)         #np.save('hw_proj0', self.projection_matrix[0])         #print("[INFO][eco.py] projection matrix[0]: \n", self.projection_matrix[0])         #print("[INFO][eco.py] projection matrix[0] shape: ", self.projection_matrix[0].shape)         self.projection_matrix = TensorList([torch.svd(C)[0][:,:cdim].clone() for C, cdim in zip(cov_x, self.compressed_dim)])                  #print("[INFO][eco.py] cov_x: \n",cov_x)                   #np.save('hw_cov_x', cov_x[0])         cov_x = x_mat @ x_mat.t()                  #print("[INFO][eco.py] x_mat2: \n",x_mat[0][0])          #np.save('hw_x_mat2', x_mat[0][0])         x_mat -= x_mat.mean(dim=1, keepdim=True)                  #print("[INFO][eco.py] x_mat mean: ", x_mat.mean(dim=1, keepdim=True)[0][0])          #print("[INFO][eco.py] x_mat1: \n",x_mat[0][0])         #np.save('hw_x_mat1', x_mat[0][0])         x_mat = TensorList([e.permute(1,0,2,3).reshape(e.shape[1], -1).clone() for e in x])         # Initialize projection matrix         #x = torch.from_numpy(x)                   #print("[INFO][eco.py] x: \n", x[0][0][0][0])         #print("[INFO][eco.py] x shape: \n", x[0].shape)         x = self.generate_init_samples(im,dpu_features)         #print("[INFO][eco.py] generate init samples")         # Extract and transform sample          self.max_scale_factor = torch.min(self.image_sz / self.base_target_sz)         self.min_scale_factor = torch.max(10 / self.base_target_sz)         self.image_sz = torch.Tensor([im.shape[2], im.shape[3]])         # Setup bounds          im = numpy_to_torch(image)         # Convert image               self.params.direction_forget_factor = (1 - max(self.params.precond_learning_rate))**self.params.CG_forgetting_rate         else:             self.params.direction_forget_factor = 0         if self.params.CG_forgetting_rate is None or max(self.params.precond_learning_rate) >= 1:         self.params.precond_learning_rate = self.fparams.attribute('learning_rate')         # Optimization options          self.yf = TensorList([dcf.label_function(sz, sig).to(self.params.device) for sz, sig in zip(self.filter_sz, sigma)])         sigma = (self.filter_sz / self.img_support_sz) * torch.sqrt(self.base_target_sz.prod()) * output_sigma_factor         output_sigma_factor = self.fparams.attribute('output_sigma_factor')         # Get label function          self.reg_energy = self.reg_filter.view(-1) @ self.reg_filter.view(-1)                                        for fparams in self.fparams])         self.reg_filter = TensorList([dcf.get_reg_filter(self.img_support_sz, self.base_target_sz, fparams).to(self.params.device) ad     q     Q       �  �  �  #  �  �  �  �  #  �  �  �  �  �  ;  �  i  J  I  -    o  n  R  0  �
  �
  �
  c
  �	  |	  �  �  �  W  V    �  e  %  $    �  �    �  k  j  5  �  �  �  �  �  u  Z  �  �  �  {  E  D  C  �  �  �  �  �  �  c  b  J  '      �  �  �  �  r  q  p                            sample_scales = self.target_scale * self.params.scale_factors         sample_pos = self.pos.round()         # Get sample          # ------- LOCALIZATION ------- #                   im = numpy_to_torch(image)         # Convert image          self.debug_info['frame_num'] = self.frame_num         self.frame_num += 1          self.debug_info = {}          track_start = time.perf_counter()     def track(self, dpu_features, image, info: dict = None) -> dict:           return out, self.img_sample_sz, sample_scales         sample_scales = self.target_scale * self.params.scale_factors         out = {'target_bbox': new_state.tolist()}          new_state = torch.cat((self.pos[[1,0]] - (self.target_sz[[1,0]]-1)/2, self.target_sz[[1,0]]))         # Return new state         self.symmetrize_filter()          self.filter_optimizer.run(self.params.post_init_CG_iter)         # Post optimization              self.filter_optimizer.run(self.params.init_CG_iter)         if not self.params.update_projection_matrix:          self.filter_optimizer.residuals = self.joint_optimizer.residuals.clone()         self.filter_optimizer.sample_energy = self.joint_problem.sample_energy         self.filter_optimizer.register(self.filter, self.training_samples, self.yf, self.sample_weights, self.reg_filter)         self.filter_optimizer = FilterOptim(self.params, self.reg_energy)         #print("[INFO][eco.py] initialize optimizer")         # Initialize optimizer              train_samp[:,:,:init_samp.shape[2],:,:] = init_samp         for train_samp, init_samp in zip(self.training_samples, compressed_samples):         compressed_samples = complex.mtimes(self.init_training_samples, self.projection_matrix)         # Re-project samples with the new projection matrix              self.joint_optimizer.run(self.params.init_CG_iter // self.params.init_GN_iter, self.params.init_GN_iter)         if self.params.update_projection_matrix:          self.joint_optimizer = GaussNewtonCG(self.joint_problem, joint_var, debug=(self.params.debug>=1), visdom=self.visdom)         joint_var = self.filter.concat(self.projection_matrix)         self.joint_problem = FactorizedConvProblem(self.init_training_samples, self.yf, self.reg_filter, self.projection_matrix, self.params, self.init_sample_weights)         #print("[INFO][eco.py] do joint optimization")         # Do joint optimization              [xf.new_zeros(1, cdim, xf.shape[2], xf.shape[3], 2) for xf, cdim in zip(train_xf, self.compressed_dim)])         self.filter = TensorList(         # Initialize filter              [xf.new_zeros(xf.shape[2], xf.shape[3], self.params.sample_memory_size, cdim, 2) for xf, cdim in zip(train_xf, self.compressed_dim)])         self.training_samples = TensorList(         # Initialize memory              sw[:num] = init_sw         for sw, init_sw, num in zip(self.sample_weights, self.init_sample_weights, num_init_samples):         self.sample_weights = TensorList([xf.new_zeros(self.params.sample_memory_size) for xf in train_xf])         self.previous_replace_ind = [None]*len(self.num_stored_samples)         self.num_stored_samples = num_init_samples         # Sample counters and weights           self.init_training_samples = train_xf.permute(2, 3, 0, 1, 4)         self.init_sample_weights = TensorList([xf.new_ones(1) / xf.shape[0] for xf in train_xf])         num_init_samples = train_xf.size(0)         # Initialize first-frame training samples          train_xf = fourier.shift_fs(train_xf, shift=shift_samp)         shift_samp = 2*math.pi * (self.pos - self.pos.round()) / (self.target_scale * self.img_support_sz)         # Shift sample                      xf[1+i:2+i,...] = fourier.shift_fs(xf[1+i:2+i,...], shift=shift_samp) 